library verilog;
use verilog.vl_types.all;
entity TestVerilog is
    port(
        first_red_pos_x : in     vl_logic_vector(9 downto 0);
        sec_red_pos_x   : in     vl_logic_vector(9 downto 0);
        top_grid_x0     : out    vl_logic_vector(9 downto 0);
        top_grid_x1     : out    vl_logic_vector(9 downto 0);
        top_grid_x2     : out    vl_logic_vector(9 downto 0);
        top_grid_x3     : out    vl_logic_vector(9 downto 0);
        top_grid_x4     : out    vl_logic_vector(9 downto 0);
        top_grid_x5     : out    vl_logic_vector(9 downto 0);
        top_grid_x6     : out    vl_logic_vector(9 downto 0);
        top_grid_x7     : out    vl_logic_vector(9 downto 0);
        top_grid_x8     : out    vl_logic_vector(9 downto 0);
        top_grid_x9     : out    vl_logic_vector(9 downto 0);
        top_grid_x10    : out    vl_logic_vector(9 downto 0);
        top_grid_x11    : out    vl_logic_vector(9 downto 0);
        top_grid_x12    : out    vl_logic_vector(9 downto 0);
        top_grid_x13    : out    vl_logic_vector(9 downto 0);
        top_grid_x14    : out    vl_logic_vector(9 downto 0);
        top_grid_x15    : out    vl_logic_vector(9 downto 0);
        top_grid_x16    : out    vl_logic_vector(9 downto 0);
        top_grid_x17    : out    vl_logic_vector(9 downto 0);
        top_grid_x18    : out    vl_logic_vector(9 downto 0);
        top_grid_x19    : out    vl_logic_vector(9 downto 0);
        top_grid_x20    : out    vl_logic_vector(9 downto 0);
        top_grid_x21    : out    vl_logic_vector(9 downto 0);
        top_grid_x22    : out    vl_logic_vector(9 downto 0);
        top_grid_x23    : out    vl_logic_vector(9 downto 0);
        top_grid_x24    : out    vl_logic_vector(9 downto 0);
        top_grid_x25    : out    vl_logic_vector(9 downto 0);
        top_grid_x26    : out    vl_logic_vector(9 downto 0);
        top_grid_x27    : out    vl_logic_vector(9 downto 0);
        top_grid_x28    : out    vl_logic_vector(9 downto 0);
        top_grid_x29    : out    vl_logic_vector(9 downto 0);
        top_grid_x30    : out    vl_logic_vector(9 downto 0);
        top_grid_x31    : out    vl_logic_vector(9 downto 0)
    );
end TestVerilog;
