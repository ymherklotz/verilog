library verilog;
use verilog.vl_types.all;
entity TestVerilog_vlg_check_tst is
    port(
        top_grid_x0     : in     vl_logic_vector(9 downto 0);
        top_grid_x1     : in     vl_logic_vector(9 downto 0);
        top_grid_x2     : in     vl_logic_vector(9 downto 0);
        top_grid_x3     : in     vl_logic_vector(9 downto 0);
        top_grid_x4     : in     vl_logic_vector(9 downto 0);
        top_grid_x5     : in     vl_logic_vector(9 downto 0);
        top_grid_x6     : in     vl_logic_vector(9 downto 0);
        top_grid_x7     : in     vl_logic_vector(9 downto 0);
        top_grid_x8     : in     vl_logic_vector(9 downto 0);
        top_grid_x9     : in     vl_logic_vector(9 downto 0);
        top_grid_x10    : in     vl_logic_vector(9 downto 0);
        top_grid_x11    : in     vl_logic_vector(9 downto 0);
        top_grid_x12    : in     vl_logic_vector(9 downto 0);
        top_grid_x13    : in     vl_logic_vector(9 downto 0);
        top_grid_x14    : in     vl_logic_vector(9 downto 0);
        top_grid_x15    : in     vl_logic_vector(9 downto 0);
        top_grid_x16    : in     vl_logic_vector(9 downto 0);
        top_grid_x17    : in     vl_logic_vector(9 downto 0);
        top_grid_x18    : in     vl_logic_vector(9 downto 0);
        top_grid_x19    : in     vl_logic_vector(9 downto 0);
        top_grid_x20    : in     vl_logic_vector(9 downto 0);
        top_grid_x21    : in     vl_logic_vector(9 downto 0);
        top_grid_x22    : in     vl_logic_vector(9 downto 0);
        top_grid_x23    : in     vl_logic_vector(9 downto 0);
        top_grid_x24    : in     vl_logic_vector(9 downto 0);
        top_grid_x25    : in     vl_logic_vector(9 downto 0);
        top_grid_x26    : in     vl_logic_vector(9 downto 0);
        top_grid_x27    : in     vl_logic_vector(9 downto 0);
        top_grid_x28    : in     vl_logic_vector(9 downto 0);
        top_grid_x29    : in     vl_logic_vector(9 downto 0);
        top_grid_x30    : in     vl_logic_vector(9 downto 0);
        top_grid_x31    : in     vl_logic_vector(9 downto 0);
        sampler_rx      : in     vl_logic
    );
end TestVerilog_vlg_check_tst;
