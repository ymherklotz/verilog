library verilog;
use verilog.vl_types.all;
entity TestVerilog_vlg_vec_tst is
end TestVerilog_vlg_vec_tst;
