// First Verilog HelloWorld Program

module hello_world;
   initial begin
	  $display("Hello World!");
	  $finish;
   end
endmodule
